`timescale 1ns / 1ps

module SectorProcessor(
  input 	clk,
  input 	reset,
// For PR		       
  input 	en_proc,
  input [2:0] 	bx_in_ProjectionRouter,
  input [59:0] 	TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout,
  input [59:0] 	TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout,
  input [7:0] 	TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout,
  input [7:0] 	TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout,
  output    TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr,
  output     TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb,
  output [7:0] TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr,
  output 	AP_L3PHIC_dataarray_data_V_wea,
  output [9:0] 	AP_L3PHIC_dataarray_data_V_writeaddr,
  output [59:0] AP_L3PHIC_dataarray_data_V_din,
  output 	AP_L3PHIC_nentries_0_V_we,
  output [7:0] 	AP_L3PHIC_nentries_0_V_din,
  output 	AP_L3PHIC_nentries_1_V_we,
  output [7:0] 	AP_L3PHIC_nentries_1_V_din,
  output 	AP_L3PHIC_nentries_2_V_we,
  output [7:0] 	AP_L3PHIC_nentries_2_V_din,
  output 	AP_L3PHIC_nentries_3_V_we,
  output [7:0] 	AP_L3PHIC_nentries_3_V_din,
  output 	AP_L3PHIC_nentries_4_V_we,
  output [7:0] 	AP_L3PHIC_nentries_4_V_din,
  output 	AP_L3PHIC_nentries_5_V_we,
  output [7:0] 	AP_L3PHIC_nentries_5_V_din,
  output 	AP_L3PHIC_nentries_6_V_we,
  output [7:0] 	AP_L3PHIC_nentries_6_V_din,
  output 	AP_L3PHIC_nentries_7_V_we,
  output [7:0] 	AP_L3PHIC_nentries_7_V_din,
// For ME
  input 	VMSME_L3PHIC17to24n1_dataarray_data_V_enb [7:0],
  input [8:0] 	VMSME_L3PHIC17to24n1_dataarray_data_V_readaddr [7:0],
  input [13:0] 	VMSME_L3PHIC17to24n1_dataarray_data_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_0_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_1_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_2_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_3_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_4_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_5_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_6_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_0_7_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_0_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_1_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_2_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_3_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_4_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_5_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_6_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_1_7_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_0_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_1_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_2_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_3_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_4_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_5_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_6_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_2_7_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_0_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_1_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_2_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_3_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_4_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_5_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_6_V_dout [7:0],
  input [3:0] 	VMSME_L3PHIC17to24n1_nentries_3_7_V_dout [7:0],
  output [2:0] 	bx_out_MatchEngine [7:0],
  output 		CM_L3PHIC17to24_dataarray_data_V_wea [7:0],
  output [7:0] 	CM_L3PHIC17to24_dataarray_data_V_writeaddr [7:0],
  output [13:0] 	CM_L3PHIC17to24_dataarray_data_V_din [7:0],
  output 		CM_L3PHIC17to24_nentries_0_V_we [7:0],
  output [6:0] 	CM_L3PHIC17to24_nentries_0_V_din [7:0],
  output 		CM_L3PHIC17to24_nentries_1_V_we [7:0],
  output [6:0] 	CM_L3PHIC17to24_nentries_1_V_din [7:0],
  output 		MatchEngine_done [7:0]		       
		     
);

//PR output
   
//wire [0:7] y2 [3:0]          // y is an 8-bit vector net with a depth of 4

  wire[2:0] bx_out_ProjectionRouter;
  reg VMPROJ_L3PHIC17to24_dataarray_data_V_wea [7:0]; //8 nonants
  wire[7:0] VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr [7:0];
  wire[20:0] VMPROJ_L3PHIC17to24_dataarray_data_V_din [7:0];
  reg VMPROJ_L3PHIC17to24_nentries_0_V_we [7:0];
  wire[7:0] VMPROJ_L3PHIC17to24_nentries_0_V_din [7:0];
  reg VMPROJ_L3PHIC17to24_nentries_1_V_we [7:0];
  wire[7:0] VMPROJ_L3PHIC17to24_nentries_1_V_din [7:0];
  reg ProjectionRouter_done;

   
ProjectionRouter_BARRELPS_BARREL_8_3_0 PR_L3PHIC(
  .ap_clk(clk),
  .ap_rst(reset),
  .ap_start(en_proc),
  .ap_done(ProjectionRouter_done),
  .bx_V(bx_in_ProjectionRouter),
  .proj1in_dataarray_data_V_ce0(TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_enb),
  .proj1in_dataarray_data_V_address0(TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_readaddr),
  .proj1in_dataarray_data_V_q0(TPROJ_L1L2XXF_L3PHIC_dataarray_data_V_dout),
  .proj1in_nentries_0_V(TPROJ_L1L2XXF_L3PHIC_nentries_0_V_dout),
  .proj1in_nentries_1_V(TPROJ_L1L2XXF_L3PHIC_nentries_1_V_dout),
  .proj2in_dataarray_data_V_ce0(TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_enb),
  .proj2in_dataarray_data_V_address0(TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_readaddr),
  .proj2in_dataarray_data_V_q0(TPROJ_L1L2XXG_L3PHIC_dataarray_data_V_dout),
  .proj2in_nentries_0_V(TPROJ_L1L2XXG_L3PHIC_nentries_0_V_dout),
  .proj2in_nentries_1_V(TPROJ_L1L2XXG_L3PHIC_nentries_1_V_dout),
  .proj3in_dataarray_data_V_ce0(TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_enb),
  .proj3in_dataarray_data_V_address0(TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_readaddr),
  .proj3in_dataarray_data_V_q0(TPROJ_L1L2XXH_L3PHIC_dataarray_data_V_dout),
  .proj3in_nentries_0_V(TPROJ_L1L2XXH_L3PHIC_nentries_0_V_dout),
  .proj3in_nentries_1_V(TPROJ_L1L2XXH_L3PHIC_nentries_1_V_dout),
  .proj4in_dataarray_data_V_ce0(TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_enb),
  .proj4in_dataarray_data_V_address0(TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_readaddr),
  .proj4in_dataarray_data_V_q0(TPROJ_L1L2XXI_L3PHIC_dataarray_data_V_dout),
  .proj4in_nentries_0_V(TPROJ_L1L2XXI_L3PHIC_nentries_0_V_dout),
  .proj4in_nentries_1_V(TPROJ_L1L2XXI_L3PHIC_nentries_1_V_dout),
  .proj5in_dataarray_data_V_ce0(TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_enb),
  .proj5in_dataarray_data_V_address0(TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_readaddr),
  .proj5in_dataarray_data_V_q0(TPROJ_L1L2XXJ_L3PHIC_dataarray_data_V_dout),
  .proj5in_nentries_0_V(TPROJ_L1L2XXJ_L3PHIC_nentries_0_V_dout),
  .proj5in_nentries_1_V(TPROJ_L1L2XXJ_L3PHIC_nentries_1_V_dout),
  .proj6in_dataarray_data_V_ce0(TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_enb),
  .proj6in_dataarray_data_V_address0(TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_readaddr),
  .proj6in_dataarray_data_V_q0(TPROJ_L5L6XXB_L3PHIC_dataarray_data_V_dout),
  .proj6in_nentries_0_V(TPROJ_L5L6XXB_L3PHIC_nentries_0_V_dout),
  .proj6in_nentries_1_V(TPROJ_L5L6XXB_L3PHIC_nentries_1_V_dout),
  .proj7in_dataarray_data_V_ce0(TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_enb),
  .proj7in_dataarray_data_V_address0(TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_readaddr),
  .proj7in_dataarray_data_V_q0(TPROJ_L5L6XXC_L3PHIC_dataarray_data_V_dout),
  .proj7in_nentries_0_V(TPROJ_L5L6XXC_L3PHIC_nentries_0_V_dout),
  .proj7in_nentries_1_V(TPROJ_L5L6XXC_L3PHIC_nentries_1_V_dout),
  .proj8in_dataarray_data_V_ce0(TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_enb),
  .proj8in_dataarray_data_V_address0(TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_readaddr),
  .proj8in_dataarray_data_V_q0(TPROJ_L5L6XXD_L3PHIC_dataarray_data_V_dout),
  .proj8in_nentries_0_V(TPROJ_L5L6XXD_L3PHIC_nentries_0_V_dout),
  .proj8in_nentries_1_V(TPROJ_L5L6XXD_L3PHIC_nentries_1_V_dout),
  .bx_o_V(bx_out_ProjectionRouter),
  .allprojout_dataarray_data_V_we0(AP_L3PHIC_dataarray_data_V_wea),
  .allprojout_dataarray_data_V_address0(AP_L3PHIC_dataarray_data_V_writeaddr),
  .allprojout_dataarray_data_V_d0(AP_L3PHIC_dataarray_data_V_din),
  .allprojout_nentries_0_V_ap_vld(AP_L3PHIC_nentries_0_V_we),
  .allprojout_nentries_0_V(AP_L3PHIC_nentries_0_V_din),
  .allprojout_nentries_1_V_ap_vld(AP_L3PHIC_nentries_1_V_we),
  .allprojout_nentries_1_V(AP_L3PHIC_nentries_1_V_din),
  .allprojout_nentries_2_V_ap_vld(AP_L3PHIC_nentries_2_V_we),
  .allprojout_nentries_2_V(AP_L3PHIC_nentries_2_V_din),
  .allprojout_nentries_3_V_ap_vld(AP_L3PHIC_nentries_3_V_we),
  .allprojout_nentries_3_V(AP_L3PHIC_nentries_3_V_din),
  .allprojout_nentries_4_V_ap_vld(AP_L3PHIC_nentries_4_V_we),
  .allprojout_nentries_4_V(AP_L3PHIC_nentries_4_V_din),
  .allprojout_nentries_5_V_ap_vld(AP_L3PHIC_nentries_5_V_we),
  .allprojout_nentries_5_V(AP_L3PHIC_nentries_5_V_din),
  .allprojout_nentries_6_V_ap_vld(AP_L3PHIC_nentries_6_V_we),
  .allprojout_nentries_6_V(AP_L3PHIC_nentries_6_V_din),
  .allprojout_nentries_7_V_ap_vld(AP_L3PHIC_nentries_7_V_we),
  .allprojout_nentries_7_V(AP_L3PHIC_nentries_7_V_din),
  .vmprojout1_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[0]),
  .vmprojout1_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[0]),
  .vmprojout1_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[0]),
  .vmprojout1_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[0]),
  .vmprojout1_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[0]),
  .vmprojout1_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[0]),
  .vmprojout1_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[0]),
  .vmprojout2_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[1]),
  .vmprojout2_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[1]),
  .vmprojout2_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[1]),
  .vmprojout2_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[1]),
  .vmprojout2_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[1]),
  .vmprojout2_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[1]),
  .vmprojout2_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[1]),
  .vmprojout3_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[2]),
  .vmprojout3_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[2]),
  .vmprojout3_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[2]),
  .vmprojout3_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[2]),
  .vmprojout3_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[2]),
  .vmprojout3_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[2]),
  .vmprojout3_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[2]),
  .vmprojout4_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[3]),
  .vmprojout4_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[3]),
  .vmprojout4_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[3]),
  .vmprojout4_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[3]),
  .vmprojout4_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[3]),
  .vmprojout4_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[3]),
  .vmprojout4_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[3]),
  .vmprojout5_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[4]),
  .vmprojout5_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[4]),
  .vmprojout5_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[4]),
  .vmprojout5_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[4]),
  .vmprojout5_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[4]),
  .vmprojout5_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[4]),
  .vmprojout5_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[4]),
  .vmprojout6_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[5]),
  .vmprojout6_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[5]),
  .vmprojout6_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[5]),
  .vmprojout6_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[5]),
  .vmprojout6_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[5]),
  .vmprojout6_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[5]),
  .vmprojout6_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[5]),
  .vmprojout7_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[6]),
  .vmprojout7_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[6]),
  .vmprojout7_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[6]),
  .vmprojout7_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[6]),
  .vmprojout7_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[6]),
  .vmprojout7_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[6]),
  .vmprojout7_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[6]),
  .vmprojout8_dataarray_data_V_we0(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[7]),
  .vmprojout8_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[7]),
  .vmprojout8_dataarray_data_V_d0(VMPROJ_L3PHIC17to24_dataarray_data_V_din[7]),
  .vmprojout8_nentries_0_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_0_V_we[7]),
  .vmprojout8_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_din[7]),
  .vmprojout8_nentries_1_V_ap_vld(VMPROJ_L3PHIC17to24_nentries_1_V_we[7]),
  .vmprojout8_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_din[7])
);


// ME Input 8 MEs
   wire VMPROJ_L3PHIC17to24_dataarray_data_V_enb [7:0];
   wire [7:0] VMPROJ_L3PHIC17to24_dataarray_data_V_readaddr [7:0];
   wire [20:0] VMPROJ_L3PHIC17to24_dataarray_data_V_dout [7:0];
   wire [6:0]  VMPROJ_L3PHIC17to24_nentries_0_V_dout [7:0];
   wire [6:0]  VMPROJ_L3PHIC17to24_nentries_1_V_dout [7:0];
   
genvar i;
   generate
      for (i=0; i<=7; i=i+1)
        begin : gen_MemoryVMProj
   Memory #(.RAM_WIDTH(21),
	    .RAM_DEPTH(256),
	    .RAM_PERFORMANCE("LOW_LATENCY"),
	    .HEX(0),
	    .INIT_FILE("")
	    ) VMPROJ_L3PHIC17to24 (
	     .clka(clk),
        .clkb(clk),
        .wea(VMPROJ_L3PHIC17to24_dataarray_data_V_wea[i]),
        .addra(VMPROJ_L3PHIC17to24_dataarray_data_V_writeaddr[i]),
        .dina(VMPROJ_L3PHIC17to24_dataarray_data_V_din[i]),
        .nent_we0(VMPROJ_L3PHIC17to24_nentries_0_V_we[i]),
        .nent_i0(VMPROJ_L3PHIC17to24_nentries_0_V_din[i]),
        .nent_we1(VMPROJ_L3PHIC17to24_nentries_1_V_we[i]),
        .nent_i1(VMPROJ_L3PHIC17to24_nentries_1_V_din[i]),
        .enb(VMPROJ_L3PHIC17to24_dataarray_data_V_enb[i]),
        .addrb(VMPROJ_L3PHIC17to24_dataarray_data_V_readaddr[i]),
        .doutb(VMPROJ_L3PHIC17to24_dataarray_data_V_dout[i]),
        .nent_o0(VMPROJ_L3PHIC17to24_nentries_0_V_dout[i]),
        .nent_o1(VMPROJ_L3PHIC17to24_nentries_1_V_dout[i]),
        .regceb(1'b1)
);
end
endgenerate   
   
  
genvar a;
generate
   for (a=0; a<=7; a=a+1)
     begin : gen_MatchEngineTopL3  
MatchEngineTopL3 MatchEngineTopL3_0( //L1 and L3 are identical, maybe should name BARRELPS
  .ap_clk(clk),
  .ap_rst(reset),
  .ap_start(ProjectionRouter_done),
  .ap_done(MatchEngine_done[a]),
  .bx_V(bx_out_ProjectionRouter),
  .bx_o_V(bx_out_MatchEngine[a]),
  .instubdata_dataarray_data_V_ce0(VMSME_L3PHIC17to24n1_dataarray_data_V_enb[a]),
  .instubdata_dataarray_data_V_address0(VMSME_L3PHIC17to24n1_dataarray_data_V_readaddr[a]),
  .instubdata_dataarray_data_V_q0(VMSME_L3PHIC17to24n1_dataarray_data_V_dout[a]),
  .instubdata_nentries_0_V_0(VMSME_L3PHIC17to24n1_nentries_0_0_V_dout[a]),
  .instubdata_nentries_0_V_1(VMSME_L3PHIC17to24n1_nentries_0_1_V_dout[a]),
  .instubdata_nentries_0_V_2(VMSME_L3PHIC17to24n1_nentries_0_2_V_dout[a]),
  .instubdata_nentries_0_V_3(VMSME_L3PHIC17to24n1_nentries_0_3_V_dout[a]),
  .instubdata_nentries_0_V_4(VMSME_L3PHIC17to24n1_nentries_0_4_V_dout[a]),
  .instubdata_nentries_0_V_5(VMSME_L3PHIC17to24n1_nentries_0_5_V_dout[a]),
  .instubdata_nentries_0_V_6(VMSME_L3PHIC17to24n1_nentries_0_6_V_dout[a]),
  .instubdata_nentries_0_V_7(VMSME_L3PHIC17to24n1_nentries_0_7_V_dout[a]),
  .instubdata_nentries_1_V_0(VMSME_L3PHIC17to24n1_nentries_1_0_V_dout[a]),
  .instubdata_nentries_1_V_1(VMSME_L3PHIC17to24n1_nentries_1_1_V_dout[a]),
  .instubdata_nentries_1_V_2(VMSME_L3PHIC17to24n1_nentries_1_2_V_dout[a]),
  .instubdata_nentries_1_V_3(VMSME_L3PHIC17to24n1_nentries_1_3_V_dout[a]),
  .instubdata_nentries_1_V_4(VMSME_L3PHIC17to24n1_nentries_1_4_V_dout[a]),
  .instubdata_nentries_1_V_5(VMSME_L3PHIC17to24n1_nentries_1_5_V_dout[a]),
  .instubdata_nentries_1_V_6(VMSME_L3PHIC17to24n1_nentries_1_6_V_dout[a]),
  .instubdata_nentries_1_V_7(VMSME_L3PHIC17to24n1_nentries_1_7_V_dout[a]),
  .instubdata_nentries_2_V_0(VMSME_L3PHIC17to24n1_nentries_2_0_V_dout[a]),
  .instubdata_nentries_2_V_1(VMSME_L3PHIC17to24n1_nentries_2_1_V_dout[a]),
  .instubdata_nentries_2_V_2(VMSME_L3PHIC17to24n1_nentries_2_2_V_dout[a]),
  .instubdata_nentries_2_V_3(VMSME_L3PHIC17to24n1_nentries_2_3_V_dout[a]),
  .instubdata_nentries_2_V_4(VMSME_L3PHIC17to24n1_nentries_2_4_V_dout[a]),
  .instubdata_nentries_2_V_5(VMSME_L3PHIC17to24n1_nentries_2_5_V_dout[a]),
  .instubdata_nentries_2_V_6(VMSME_L3PHIC17to24n1_nentries_2_6_V_dout[a]),
  .instubdata_nentries_2_V_7(VMSME_L3PHIC17to24n1_nentries_2_7_V_dout[a]),
  .instubdata_nentries_3_V_0(VMSME_L3PHIC17to24n1_nentries_3_0_V_dout[a]),
  .instubdata_nentries_3_V_1(VMSME_L3PHIC17to24n1_nentries_3_1_V_dout[a]),
  .instubdata_nentries_3_V_2(VMSME_L3PHIC17to24n1_nentries_3_2_V_dout[a]),
  .instubdata_nentries_3_V_3(VMSME_L3PHIC17to24n1_nentries_3_3_V_dout[a]),
  .instubdata_nentries_3_V_4(VMSME_L3PHIC17to24n1_nentries_3_4_V_dout[a]),
  .instubdata_nentries_3_V_5(VMSME_L3PHIC17to24n1_nentries_3_5_V_dout[a]),
  .instubdata_nentries_3_V_6(VMSME_L3PHIC17to24n1_nentries_3_6_V_dout[a]),
  .instubdata_nentries_3_V_7(VMSME_L3PHIC17to24n1_nentries_3_7_V_dout[a]),				      
  .inprojdata_dataarray_data_V_ce0(VMPROJ_L3PHIC17to24_dataarray_data_V_enb[a]),
  .inprojdata_dataarray_data_V_address0(VMPROJ_L3PHIC17to24_dataarray_data_V_readaddr[a]),
  .inprojdata_dataarray_data_V_q0(VMPROJ_L3PHIC17to24_dataarray_data_V_dout[a]),
  .inprojdata_nentries_0_V(VMPROJ_L3PHIC17to24_nentries_0_V_dout[a]),
  .inprojdata_nentries_1_V(VMPROJ_L3PHIC17to24_nentries_1_V_dout[a]),
  .outcandmatch_dataarray_data_V_we0(CM_L3PHIC17to24_dataarray_data_V_wea[a]),
  .outcandmatch_dataarray_data_V_address0(CM_L3PHIC17to24_dataarray_data_V_writeaddr[a]),
  .outcandmatch_dataarray_data_V_d0(CM_L3PHIC17to24_dataarray_data_V_din[a]),
  .outcandmatch_nentries_0_V_ap_vld(CM_L3PHIC17to24_nentries_0_V_we[a]),
  .outcandmatch_nentries_0_V(CM_L3PHIC17to24_nentries_0_V_din[a]),
  .outcandmatch_nentries_1_V_ap_vld(CM_L3PHIC17to24_nentries_1_V_we[a]),
  .outcandmatch_nentries_1_V(CM_L3PHIC17to24_nentries_1_V_din[a])
);
end
endgenerate

endmodule
