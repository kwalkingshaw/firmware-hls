`timescale 1ns / 1ps

module SectorProcessor(
  input 	clk,
  input 	reset,
  input 	en_proc,
  input [2:0] 	bx_in_MatchEngine,
  output 	VMSME_L1PHIE20n1_dataarray_data_V_enb,
  output [8:0] 	VMSME_L1PHIE20n1_dataarray_data_V_readaddr,
  input [13:0] 	VMSME_L1PHIE20n1_dataarray_data_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_0_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_1_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_2_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_3_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_4_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_5_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_6_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_0_7_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_0_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_1_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_2_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_3_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_4_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_5_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_6_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_1_7_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_0_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_1_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_2_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_3_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_4_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_5_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_6_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_2_7_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_0_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_1_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_2_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_3_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_4_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_5_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_6_V_dout,
  input [3:0] 	VMSME_L1PHIE20n1_nentries_3_7_V_dout,
  output 	VMPROJ_L1PHIE20_dataarray_data_V_enb,
  output [7:0] 	VMPROJ_L1PHIE20_dataarray_data_V_readaddr,
  input [20:0] 	VMPROJ_L1PHIE20_dataarray_data_V_dout,
  input [6:0] 	VMPROJ_L1PHIE20_nentries_0_V_dout,
  input [6:0] 	VMPROJ_L1PHIE20_nentries_1_V_dout,
  output [2:0] 	bx_out_MatchEngine,
  output 	CM_L1PHIE20_dataarray_data_V_wea,
  output [7:0] 	CM_L1PHIE20_dataarray_data_V_writeaddr,
  output [13:0] CM_L1PHIE20_dataarray_data_V_din,
  output 	CM_L1PHIE20_nentries_0_V_we,
  output [6:0] 	CM_L1PHIE20_nentries_0_V_din,
  output 	CM_L1PHIE20_nentries_1_V_we,
  output [6:0] 	CM_L1PHIE20_nentries_1_V_din,
  output 	MatchEngine_done
);

MatchEngineTopL1_0 MatchEngineTopL1_0(
  .ap_clk(clk),
  .ap_rst(reset),
  .ap_start(en_proc),
  .ap_done(MatchEngine_done),
  .bx_V(bx_in_MatchEngine),
  .bx_o_V(bx_out_MatchEngine),
  .instubdata_dataarray_data_V_ce0(VMSME_L1PHIE20n1_dataarray_data_V_enb),
  .instubdata_dataarray_data_V_address0(VMSME_L1PHIE20n1_dataarray_data_V_readaddr),
  .instubdata_dataarray_data_V_q0(VMSME_L1PHIE20n1_dataarray_data_V_dout),
  .instubdata_nentries_0_V_0(VMSME_L1PHIE20n1_nentries_0_0_V_dout),
  .instubdata_nentries_0_V_1(VMSME_L1PHIE20n1_nentries_0_1_V_dout),
  .instubdata_nentries_0_V_2(VMSME_L1PHIE20n1_nentries_0_2_V_dout),
  .instubdata_nentries_0_V_3(VMSME_L1PHIE20n1_nentries_0_3_V_dout),
  .instubdata_nentries_0_V_4(VMSME_L1PHIE20n1_nentries_0_4_V_dout),
  .instubdata_nentries_0_V_5(VMSME_L1PHIE20n1_nentries_0_5_V_dout),
  .instubdata_nentries_0_V_6(VMSME_L1PHIE20n1_nentries_0_6_V_dout),
  .instubdata_nentries_0_V_7(VMSME_L1PHIE20n1_nentries_0_7_V_dout),
  .instubdata_nentries_1_V_0(VMSME_L1PHIE20n1_nentries_1_0_V_dout),
  .instubdata_nentries_1_V_1(VMSME_L1PHIE20n1_nentries_1_1_V_dout),
  .instubdata_nentries_1_V_2(VMSME_L1PHIE20n1_nentries_1_2_V_dout),
  .instubdata_nentries_1_V_3(VMSME_L1PHIE20n1_nentries_1_3_V_dout),
  .instubdata_nentries_1_V_4(VMSME_L1PHIE20n1_nentries_1_4_V_dout),
  .instubdata_nentries_1_V_5(VMSME_L1PHIE20n1_nentries_1_5_V_dout),
  .instubdata_nentries_1_V_6(VMSME_L1PHIE20n1_nentries_1_6_V_dout),
  .instubdata_nentries_1_V_7(VMSME_L1PHIE20n1_nentries_1_7_V_dout),
  .instubdata_nentries_2_V_0(VMSME_L1PHIE20n1_nentries_2_0_V_dout),
  .instubdata_nentries_2_V_1(VMSME_L1PHIE20n1_nentries_2_1_V_dout),
  .instubdata_nentries_2_V_2(VMSME_L1PHIE20n1_nentries_2_2_V_dout),
  .instubdata_nentries_2_V_3(VMSME_L1PHIE20n1_nentries_2_3_V_dout),
  .instubdata_nentries_2_V_4(VMSME_L1PHIE20n1_nentries_2_4_V_dout),
  .instubdata_nentries_2_V_5(VMSME_L1PHIE20n1_nentries_2_5_V_dout),
  .instubdata_nentries_2_V_6(VMSME_L1PHIE20n1_nentries_2_6_V_dout),
  .instubdata_nentries_2_V_7(VMSME_L1PHIE20n1_nentries_2_7_V_dout),
  .instubdata_nentries_3_V_0(VMSME_L1PHIE20n1_nentries_3_0_V_dout),
  .instubdata_nentries_3_V_1(VMSME_L1PHIE20n1_nentries_3_1_V_dout),
  .instubdata_nentries_3_V_2(VMSME_L1PHIE20n1_nentries_3_2_V_dout),
  .instubdata_nentries_3_V_3(VMSME_L1PHIE20n1_nentries_3_3_V_dout),
  .instubdata_nentries_3_V_4(VMSME_L1PHIE20n1_nentries_3_4_V_dout),
  .instubdata_nentries_3_V_5(VMSME_L1PHIE20n1_nentries_3_5_V_dout),
  .instubdata_nentries_3_V_6(VMSME_L1PHIE20n1_nentries_3_6_V_dout),
  .instubdata_nentries_3_V_7(VMSME_L1PHIE20n1_nentries_3_7_V_dout),				      
  .inprojdata_dataarray_data_V_ce0(VMPROJ_L1PHIE20_dataarray_data_V_enb),
  .inprojdata_dataarray_data_V_address0(VMPROJ_L1PHIE20_dataarray_data_V_readaddr),
  .inprojdata_dataarray_data_V_q0(VMPROJ_L1PHIE20_dataarray_data_V_dout),
  .inprojdata_nentries_0_V(VMPROJ_L1PHIE20_nentries_0_V_dout),
  .inprojdata_nentries_1_V(VMPROJ_L1PHIE20_nentries_1_V_dout),
  .outcandmatch_dataarray_data_V_we0(CM_L1PHIE20_dataarray_data_V_wea),
  .outcandmatch_dataarray_data_V_address0(CM_L1PHIE20_dataarray_data_V_writeaddr),
  .outcandmatch_dataarray_data_V_d0(CM_L1PHIE20_dataarray_data_V_din),
  .outcandmatch_nentries_0_V_ap_vld(CM_L1PHIE20_nentries_0_V_we),
  .outcandmatch_nentries_0_V(CM_L1PHIE20_nentries_0_V_din),
  .outcandmatch_nentries_1_V_ap_vld(CM_L1PHIE20_nentries_1_V_we),
  .outcandmatch_nentries_1_V(CM_L1PHIE20_nentries_1_V_din)
);

endmodule
